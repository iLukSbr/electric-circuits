* Netlist E:\Pastas\Documentos\UTFPR\4Per\Circuitos El�tricos ELEB21-S72\Listas de Exerc�cios\Atividade Complementar Bode\ativ_simu.psimsch *

.include "C:\Altair\Altair_PSIM_2023.1\SPICElib\PSIM_SPICE.sub"

.ac dec 10000 1000 8000
V_V1 1 2 SINE( 0 0.3988 1000 0 0 0 )
R_R1 1 3 40
L_L1 3 4 0.03
C_C1 4 2 1E-07

* Matching PSIM probes to SPICE probes *

.end
