* C:\Users\lucas\Desktop\p2\1.sch

* Schematics Version 9.1 - Web Update 1
* Thu Jun 27 10:22:25 2024



** Analysis setup **
.tran 10ms 30s 0 1ms


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "1.net"
.INC "1.als"


.probe


.END
